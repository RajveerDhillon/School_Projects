library verilog;
use verilog.vl_types.all;
entity lab_1f_vlg_vec_tst is
end lab_1f_vlg_vec_tst;
