library verilog;
use verilog.vl_types.all;
entity registerPC_vlg_vec_tst is
end registerPC_vlg_vec_tst;
