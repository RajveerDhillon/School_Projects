library verilog;
use verilog.vl_types.all;
entity uze_vlg_vec_tst is
end uze_vlg_vec_tst;
