library verilog;
use verilog.vl_types.all;
entity lab_1f is
    port(
        f               : out    vl_logic;
        w1              : in     vl_logic;
        w2              : in     vl_logic;
        w3              : in     vl_logic;
        w4              : in     vl_logic;
        x2              : in     vl_logic
    );
end lab_1f;
