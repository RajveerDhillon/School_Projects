library verilog;
use verilog.vl_types.all;
entity lab_one_vlg_vec_tst is
end lab_one_vlg_vec_tst;
