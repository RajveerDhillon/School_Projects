library verilog;
use verilog.vl_types.all;
entity reg1_vlg_vec_tst is
end reg1_vlg_vec_tst;
