library verilog;
use verilog.vl_types.all;
entity leftSH_vlg_vec_tst is
end leftSH_vlg_vec_tst;
