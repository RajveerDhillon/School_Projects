LIBRARY ieee ;
USE ieee.std_logic_1164.all ;
ENTITY ALUDE IS
PORT ( S: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
       Z,X : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)) ;
END ALUDE ;
ARCHITECTURE Behavior OF ALUDE IS
 BEGIN
Z<= S(3 DOWNTO 0);
X<= S(7 DOWNTO 4);
END Behavior ;