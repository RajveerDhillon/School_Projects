library verilog;
use verilog.vl_types.all;
entity rightSH_vlg_vec_tst is
end rightSH_vlg_vec_tst;
