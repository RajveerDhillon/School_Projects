library verilog;
use verilog.vl_types.all;
entity lab4Bvd_vlg_vec_tst is
end lab4Bvd_vlg_vec_tst;
