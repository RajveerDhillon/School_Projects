library verilog;
use verilog.vl_types.all;
entity testbench_vlg_vec_tst is
end testbench_vlg_vec_tst;
