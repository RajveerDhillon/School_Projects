library verilog;
use verilog.vl_types.all;
entity reducer_vlg_vec_tst is
end reducer_vlg_vec_tst;
