library verilog;
use verilog.vl_types.all;
entity and32_vlg_vec_tst is
end and32_vlg_vec_tst;
