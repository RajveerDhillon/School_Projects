library verilog;
use verilog.vl_types.all;
entity lab_1f_vlg_check_tst is
    port(
        f               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab_1f_vlg_check_tst;
