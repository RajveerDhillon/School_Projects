library verilog;
use verilog.vl_types.all;
entity lze_vlg_vec_tst is
end lze_vlg_vec_tst;
