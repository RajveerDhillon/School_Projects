library verilog;
use verilog.vl_types.all;
entity lab4b_vlg_check_tst is
    port(
        CarryOut        : in     vl_logic;
        Zero            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab4b_vlg_check_tst;
