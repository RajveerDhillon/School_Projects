
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity C is
port ( 
A, B, C, D : in std_logic;
f : OUT std_logic );
end C;
architecture Behavioral of C is

begin
process 
BEGIN 

end process;
end Behavioral;
