library verilog;
use verilog.vl_types.all;
entity lab1_first_part_vlg_vec_tst is
end lab1_first_part_vlg_vec_tst;
