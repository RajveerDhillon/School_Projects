library verilog;
use verilog.vl_types.all;
entity lab_1f_vlg_sample_tst is
    port(
        w1              : in     vl_logic;
        w2              : in     vl_logic;
        w3              : in     vl_logic;
        w4              : in     vl_logic;
        x2              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end lab_1f_vlg_sample_tst;
