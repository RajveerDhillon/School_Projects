library verilog;
use verilog.vl_types.all;
entity lab4b_vlg_vec_tst is
end lab4b_vlg_vec_tst;
