library verilog;
use verilog.vl_types.all;
entity or32_vlg_vec_tst is
end or32_vlg_vec_tst;
